library ieee;
use ieee.std_logic_1146.all;
use ieee.numeric_std.all;




